
module sum_product();

   integer a;
   integer b;
   integer sum;
   
   initial begin
   a=5;
   b=1;
   sum=a+b;
   $display("\n\t %0d + %0d =%0d",a,b,sum);
   end
endmodule

   